// Solution by Seunghyeok Lee
// Problem: If statement latches
// Problem link: https://hdlbits.01xz.net/wiki/Always_if2

module top_module (
    input      cpu_overheated,
    output reg shut_off_computer,
    input      arrived,
    input      gas_tank_empty,
    output reg keep_driving 
);

    // because we specify the else case, no latch is used
    always @(*) begin
        if (cpu_overheated)
           shut_off_computer = 1;
        else
            shut_off_computer = 0; 
    end

    always @(*) begin
        if (~arrived)
           keep_driving = ~gas_tank_empty;
        else
            keep_driving = 0;
    end

endmodule
