// Solution by Seunghyeok Lee
// Problem: Simple Wire

module top_module ( input in, output out );
    assign out = in;
endmodule